
/*
    file name  : core_pkg.sv
    Description: core_pkg contains parameters, functions
*/

package core_pkg;



endpackage
